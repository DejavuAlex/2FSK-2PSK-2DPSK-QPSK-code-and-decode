module test(
    output[7:0]a,
	 output[7:0]HEX0
	);
	assign a=2'h07;
	assign HEX0=a;
endmodule
	