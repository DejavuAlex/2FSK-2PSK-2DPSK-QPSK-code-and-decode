module seq(
    input clk,
    output seq
);







endmodule
